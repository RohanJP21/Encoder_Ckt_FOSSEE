* C:\Users\mistr\eSim-Workspace\encoder\encoder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/14/21 21:35:05

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  Net-_U4-Pad4_ Net-_U4-Pad5_ Net-_U5-Pad3_ d_or		
U6  Net-_U4-Pad4_ Net-_U4-Pad6_ Net-_U6-Pad3_ d_or		
U7  Net-_U5-Pad3_ Net-_U6-Pad3_ A1 A0 dac_bridge_2		
U4  Y3 Y2 Y1 Net-_U4-Pad4_ Net-_U4-Pad5_ Net-_U4-Pad6_ adc_bridge_3		
R1  A1 GND eSim_R		
R2  A0 GND eSim_R		
v1  Y3 GND DC		
v2  Y2 GND DC		
v3  Y1 GND DC		
U1  Y3 plot_v1		
U2  Y2 plot_v1		
U3  Y1 plot_v1		
U8  A0 plot_v1		
U9  A1 plot_v1		

.end
